module i2c (
	input reg scl,
	input reg sda
);
	reg [3:0] state;

		
endmodule

